library verilog;
use verilog.vl_types.all;
entity fp_add_sub_vlg_vec_tst is
end fp_add_sub_vlg_vec_tst;
