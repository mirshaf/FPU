library verilog;
use verilog.vl_types.all;
entity unsigned_multiplier_vlg_vec_tst is
end unsigned_multiplier_vlg_vec_tst;
