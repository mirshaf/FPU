library verilog;
use verilog.vl_types.all;
entity fp_mul_vlg_vec_tst is
end fp_mul_vlg_vec_tst;
