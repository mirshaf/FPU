library verilog;
use verilog.vl_types.all;
entity FPU_vlg_vec_tst is
end FPU_vlg_vec_tst;
